`timescale 1ns / 1ps

module NextState #(parameter map_width = 8)
    (
    input [map_width**2-1:0] state_in,
    output [map_width**2-1:0] state_out
    );
    
    function solve_cell(input [8:0] cell_state);
    begin
        case (cell_state)
            9'b000000000: solve_cell = 0;
            9'b000000001: solve_cell = 0;
            9'b000000010: solve_cell = 0;
            9'b000000011: solve_cell = 0;
            9'b000000100: solve_cell = 0;
            9'b000000101: solve_cell = 0;
            9'b000000110: solve_cell = 0;
            9'b000000111: solve_cell = 1;
            9'b000001000: solve_cell = 0;
            9'b000001001: solve_cell = 0;
            9'b000001010: solve_cell = 0;
            9'b000001011: solve_cell = 1;
            9'b000001100: solve_cell = 0;
            9'b000001101: solve_cell = 1;
            9'b000001110: solve_cell = 1;
            9'b000001111: solve_cell = 0;
            9'b000010000: solve_cell = 0;
            9'b000010001: solve_cell = 0;
            9'b000010010: solve_cell = 0;
            9'b000010011: solve_cell = 1;
            9'b000010100: solve_cell = 0;
            9'b000010101: solve_cell = 1;
            9'b000010110: solve_cell = 1;
            9'b000010111: solve_cell = 1;
            9'b000011000: solve_cell = 0;
            9'b000011001: solve_cell = 1;
            9'b000011010: solve_cell = 1;
            9'b000011011: solve_cell = 1;
            9'b000011100: solve_cell = 1;
            9'b000011101: solve_cell = 1;
            9'b000011110: solve_cell = 1;
            9'b000011111: solve_cell = 0;
            9'b000100000: solve_cell = 0;
            9'b000100001: solve_cell = 0;
            9'b000100010: solve_cell = 0;
            9'b000100011: solve_cell = 1;
            9'b000100100: solve_cell = 0;
            9'b000100101: solve_cell = 1;
            9'b000100110: solve_cell = 1;
            9'b000100111: solve_cell = 0;
            9'b000101000: solve_cell = 0;
            9'b000101001: solve_cell = 1;
            9'b000101010: solve_cell = 1;
            9'b000101011: solve_cell = 0;
            9'b000101100: solve_cell = 1;
            9'b000101101: solve_cell = 0;
            9'b000101110: solve_cell = 0;
            9'b000101111: solve_cell = 0;
            9'b000110000: solve_cell = 0;
            9'b000110001: solve_cell = 1;
            9'b000110010: solve_cell = 1;
            9'b000110011: solve_cell = 1;
            9'b000110100: solve_cell = 1;
            9'b000110101: solve_cell = 1;
            9'b000110110: solve_cell = 1;
            9'b000110111: solve_cell = 0;
            9'b000111000: solve_cell = 1;
            9'b000111001: solve_cell = 1;
            9'b000111010: solve_cell = 1;
            9'b000111011: solve_cell = 0;
            9'b000111100: solve_cell = 1;
            9'b000111101: solve_cell = 0;
            9'b000111110: solve_cell = 0;
            9'b000111111: solve_cell = 0;
            9'b001000000: solve_cell = 0;
            9'b001000001: solve_cell = 0;
            9'b001000010: solve_cell = 0;
            9'b001000011: solve_cell = 1;
            9'b001000100: solve_cell = 0;
            9'b001000101: solve_cell = 1;
            9'b001000110: solve_cell = 1;
            9'b001000111: solve_cell = 0;
            9'b001001000: solve_cell = 0;
            9'b001001001: solve_cell = 1;
            9'b001001010: solve_cell = 1;
            9'b001001011: solve_cell = 0;
            9'b001001100: solve_cell = 1;
            9'b001001101: solve_cell = 0;
            9'b001001110: solve_cell = 0;
            9'b001001111: solve_cell = 0;
            9'b001010000: solve_cell = 0;
            9'b001010001: solve_cell = 1;
            9'b001010010: solve_cell = 1;
            9'b001010011: solve_cell = 1;
            9'b001010100: solve_cell = 1;
            9'b001010101: solve_cell = 1;
            9'b001010110: solve_cell = 1;
            9'b001010111: solve_cell = 0;
            9'b001011000: solve_cell = 1;
            9'b001011001: solve_cell = 1;
            9'b001011010: solve_cell = 1;
            9'b001011011: solve_cell = 0;
            9'b001011100: solve_cell = 1;
            9'b001011101: solve_cell = 0;
            9'b001011110: solve_cell = 0;
            9'b001011111: solve_cell = 0;
            9'b001100000: solve_cell = 0;
            9'b001100001: solve_cell = 1;
            9'b001100010: solve_cell = 1;
            9'b001100011: solve_cell = 0;
            9'b001100100: solve_cell = 1;
            9'b001100101: solve_cell = 0;
            9'b001100110: solve_cell = 0;
            9'b001100111: solve_cell = 0;
            9'b001101000: solve_cell = 1;
            9'b001101001: solve_cell = 0;
            9'b001101010: solve_cell = 0;
            9'b001101011: solve_cell = 0;
            9'b001101100: solve_cell = 0;
            9'b001101101: solve_cell = 0;
            9'b001101110: solve_cell = 0;
            9'b001101111: solve_cell = 0;
            9'b001110000: solve_cell = 1;
            9'b001110001: solve_cell = 1;
            9'b001110010: solve_cell = 1;
            9'b001110011: solve_cell = 0;
            9'b001110100: solve_cell = 1;
            9'b001110101: solve_cell = 0;
            9'b001110110: solve_cell = 0;
            9'b001110111: solve_cell = 0;
            9'b001111000: solve_cell = 1;
            9'b001111001: solve_cell = 0;
            9'b001111010: solve_cell = 0;
            9'b001111011: solve_cell = 0;
            9'b001111100: solve_cell = 0;
            9'b001111101: solve_cell = 0;
            9'b001111110: solve_cell = 0;
            9'b001111111: solve_cell = 0;
            9'b010000000: solve_cell = 0;
            9'b010000001: solve_cell = 0;
            9'b010000010: solve_cell = 0;
            9'b010000011: solve_cell = 1;
            9'b010000100: solve_cell = 0;
            9'b010000101: solve_cell = 1;
            9'b010000110: solve_cell = 1;
            9'b010000111: solve_cell = 0;
            9'b010001000: solve_cell = 0;
            9'b010001001: solve_cell = 1;
            9'b010001010: solve_cell = 1;
            9'b010001011: solve_cell = 0;
            9'b010001100: solve_cell = 1;
            9'b010001101: solve_cell = 0;
            9'b010001110: solve_cell = 0;
            9'b010001111: solve_cell = 0;
            9'b010010000: solve_cell = 0;
            9'b010010001: solve_cell = 1;
            9'b010010010: solve_cell = 1;
            9'b010010011: solve_cell = 1;
            9'b010010100: solve_cell = 1;
            9'b010010101: solve_cell = 1;
            9'b010010110: solve_cell = 1;
            9'b010010111: solve_cell = 0;
            9'b010011000: solve_cell = 1;
            9'b010011001: solve_cell = 1;
            9'b010011010: solve_cell = 1;
            9'b010011011: solve_cell = 0;
            9'b010011100: solve_cell = 1;
            9'b010011101: solve_cell = 0;
            9'b010011110: solve_cell = 0;
            9'b010011111: solve_cell = 0;
            9'b010100000: solve_cell = 0;
            9'b010100001: solve_cell = 1;
            9'b010100010: solve_cell = 1;
            9'b010100011: solve_cell = 0;
            9'b010100100: solve_cell = 1;
            9'b010100101: solve_cell = 0;
            9'b010100110: solve_cell = 0;
            9'b010100111: solve_cell = 0;
            9'b010101000: solve_cell = 1;
            9'b010101001: solve_cell = 0;
            9'b010101010: solve_cell = 0;
            9'b010101011: solve_cell = 0;
            9'b010101100: solve_cell = 0;
            9'b010101101: solve_cell = 0;
            9'b010101110: solve_cell = 0;
            9'b010101111: solve_cell = 0;
            9'b010110000: solve_cell = 1;
            9'b010110001: solve_cell = 1;
            9'b010110010: solve_cell = 1;
            9'b010110011: solve_cell = 0;
            9'b010110100: solve_cell = 1;
            9'b010110101: solve_cell = 0;
            9'b010110110: solve_cell = 0;
            9'b010110111: solve_cell = 0;
            9'b010111000: solve_cell = 1;
            9'b010111001: solve_cell = 0;
            9'b010111010: solve_cell = 0;
            9'b010111011: solve_cell = 0;
            9'b010111100: solve_cell = 0;
            9'b010111101: solve_cell = 0;
            9'b010111110: solve_cell = 0;
            9'b010111111: solve_cell = 0;
            9'b011000000: solve_cell = 0;
            9'b011000001: solve_cell = 1;
            9'b011000010: solve_cell = 1;
            9'b011000011: solve_cell = 0;
            9'b011000100: solve_cell = 1;
            9'b011000101: solve_cell = 0;
            9'b011000110: solve_cell = 0;
            9'b011000111: solve_cell = 0;
            9'b011001000: solve_cell = 1;
            9'b011001001: solve_cell = 0;
            9'b011001010: solve_cell = 0;
            9'b011001011: solve_cell = 0;
            9'b011001100: solve_cell = 0;
            9'b011001101: solve_cell = 0;
            9'b011001110: solve_cell = 0;
            9'b011001111: solve_cell = 0;
            9'b011010000: solve_cell = 1;
            9'b011010001: solve_cell = 1;
            9'b011010010: solve_cell = 1;
            9'b011010011: solve_cell = 0;
            9'b011010100: solve_cell = 1;
            9'b011010101: solve_cell = 0;
            9'b011010110: solve_cell = 0;
            9'b011010111: solve_cell = 0;
            9'b011011000: solve_cell = 1;
            9'b011011001: solve_cell = 0;
            9'b011011010: solve_cell = 0;
            9'b011011011: solve_cell = 0;
            9'b011011100: solve_cell = 0;
            9'b011011101: solve_cell = 0;
            9'b011011110: solve_cell = 0;
            9'b011011111: solve_cell = 0;
            9'b011100000: solve_cell = 1;
            9'b011100001: solve_cell = 0;
            9'b011100010: solve_cell = 0;
            9'b011100011: solve_cell = 0;
            9'b011100100: solve_cell = 0;
            9'b011100101: solve_cell = 0;
            9'b011100110: solve_cell = 0;
            9'b011100111: solve_cell = 0;
            9'b011101000: solve_cell = 0;
            9'b011101001: solve_cell = 0;
            9'b011101010: solve_cell = 0;
            9'b011101011: solve_cell = 0;
            9'b011101100: solve_cell = 0;
            9'b011101101: solve_cell = 0;
            9'b011101110: solve_cell = 0;
            9'b011101111: solve_cell = 0;
            9'b011110000: solve_cell = 1;
            9'b011110001: solve_cell = 0;
            9'b011110010: solve_cell = 0;
            9'b011110011: solve_cell = 0;
            9'b011110100: solve_cell = 0;
            9'b011110101: solve_cell = 0;
            9'b011110110: solve_cell = 0;
            9'b011110111: solve_cell = 0;
            9'b011111000: solve_cell = 0;
            9'b011111001: solve_cell = 0;
            9'b011111010: solve_cell = 0;
            9'b011111011: solve_cell = 0;
            9'b011111100: solve_cell = 0;
            9'b011111101: solve_cell = 0;
            9'b011111110: solve_cell = 0;
            9'b011111111: solve_cell = 0;
            9'b100000000: solve_cell = 0;
            9'b100000001: solve_cell = 0;
            9'b100000010: solve_cell = 0;
            9'b100000011: solve_cell = 1;
            9'b100000100: solve_cell = 0;
            9'b100000101: solve_cell = 1;
            9'b100000110: solve_cell = 1;
            9'b100000111: solve_cell = 0;
            9'b100001000: solve_cell = 0;
            9'b100001001: solve_cell = 1;
            9'b100001010: solve_cell = 1;
            9'b100001011: solve_cell = 0;
            9'b100001100: solve_cell = 1;
            9'b100001101: solve_cell = 0;
            9'b100001110: solve_cell = 0;
            9'b100001111: solve_cell = 0;
            9'b100010000: solve_cell = 0;
            9'b100010001: solve_cell = 1;
            9'b100010010: solve_cell = 1;
            9'b100010011: solve_cell = 1;
            9'b100010100: solve_cell = 1;
            9'b100010101: solve_cell = 1;
            9'b100010110: solve_cell = 1;
            9'b100010111: solve_cell = 0;
            9'b100011000: solve_cell = 1;
            9'b100011001: solve_cell = 1;
            9'b100011010: solve_cell = 1;
            9'b100011011: solve_cell = 0;
            9'b100011100: solve_cell = 1;
            9'b100011101: solve_cell = 0;
            9'b100011110: solve_cell = 0;
            9'b100011111: solve_cell = 0;
            9'b100100000: solve_cell = 0;
            9'b100100001: solve_cell = 1;
            9'b100100010: solve_cell = 1;
            9'b100100011: solve_cell = 0;
            9'b100100100: solve_cell = 1;
            9'b100100101: solve_cell = 0;
            9'b100100110: solve_cell = 0;
            9'b100100111: solve_cell = 0;
            9'b100101000: solve_cell = 1;
            9'b100101001: solve_cell = 0;
            9'b100101010: solve_cell = 0;
            9'b100101011: solve_cell = 0;
            9'b100101100: solve_cell = 0;
            9'b100101101: solve_cell = 0;
            9'b100101110: solve_cell = 0;
            9'b100101111: solve_cell = 0;
            9'b100110000: solve_cell = 1;
            9'b100110001: solve_cell = 1;
            9'b100110010: solve_cell = 1;
            9'b100110011: solve_cell = 0;
            9'b100110100: solve_cell = 1;
            9'b100110101: solve_cell = 0;
            9'b100110110: solve_cell = 0;
            9'b100110111: solve_cell = 0;
            9'b100111000: solve_cell = 1;
            9'b100111001: solve_cell = 0;
            9'b100111010: solve_cell = 0;
            9'b100111011: solve_cell = 0;
            9'b100111100: solve_cell = 0;
            9'b100111101: solve_cell = 0;
            9'b100111110: solve_cell = 0;
            9'b100111111: solve_cell = 0;
            9'b101000000: solve_cell = 0;
            9'b101000001: solve_cell = 1;
            9'b101000010: solve_cell = 1;
            9'b101000011: solve_cell = 0;
            9'b101000100: solve_cell = 1;
            9'b101000101: solve_cell = 0;
            9'b101000110: solve_cell = 0;
            9'b101000111: solve_cell = 0;
            9'b101001000: solve_cell = 1;
            9'b101001001: solve_cell = 0;
            9'b101001010: solve_cell = 0;
            9'b101001011: solve_cell = 0;
            9'b101001100: solve_cell = 0;
            9'b101001101: solve_cell = 0;
            9'b101001110: solve_cell = 0;
            9'b101001111: solve_cell = 0;
            9'b101010000: solve_cell = 1;
            9'b101010001: solve_cell = 1;
            9'b101010010: solve_cell = 1;
            9'b101010011: solve_cell = 0;
            9'b101010100: solve_cell = 1;
            9'b101010101: solve_cell = 0;
            9'b101010110: solve_cell = 0;
            9'b101010111: solve_cell = 0;
            9'b101011000: solve_cell = 1;
            9'b101011001: solve_cell = 0;
            9'b101011010: solve_cell = 0;
            9'b101011011: solve_cell = 0;
            9'b101011100: solve_cell = 0;
            9'b101011101: solve_cell = 0;
            9'b101011110: solve_cell = 0;
            9'b101011111: solve_cell = 0;
            9'b101100000: solve_cell = 1;
            9'b101100001: solve_cell = 0;
            9'b101100010: solve_cell = 0;
            9'b101100011: solve_cell = 0;
            9'b101100100: solve_cell = 0;
            9'b101100101: solve_cell = 0;
            9'b101100110: solve_cell = 0;
            9'b101100111: solve_cell = 0;
            9'b101101000: solve_cell = 0;
            9'b101101001: solve_cell = 0;
            9'b101101010: solve_cell = 0;
            9'b101101011: solve_cell = 0;
            9'b101101100: solve_cell = 0;
            9'b101101101: solve_cell = 0;
            9'b101101110: solve_cell = 0;
            9'b101101111: solve_cell = 0;
            9'b101110000: solve_cell = 1;
            9'b101110001: solve_cell = 0;
            9'b101110010: solve_cell = 0;
            9'b101110011: solve_cell = 0;
            9'b101110100: solve_cell = 0;
            9'b101110101: solve_cell = 0;
            9'b101110110: solve_cell = 0;
            9'b101110111: solve_cell = 0;
            9'b101111000: solve_cell = 0;
            9'b101111001: solve_cell = 0;
            9'b101111010: solve_cell = 0;
            9'b101111011: solve_cell = 0;
            9'b101111100: solve_cell = 0;
            9'b101111101: solve_cell = 0;
            9'b101111110: solve_cell = 0;
            9'b101111111: solve_cell = 0;
            9'b110000000: solve_cell = 0;
            9'b110000001: solve_cell = 1;
            9'b110000010: solve_cell = 1;
            9'b110000011: solve_cell = 0;
            9'b110000100: solve_cell = 1;
            9'b110000101: solve_cell = 0;
            9'b110000110: solve_cell = 0;
            9'b110000111: solve_cell = 0;
            9'b110001000: solve_cell = 1;
            9'b110001001: solve_cell = 0;
            9'b110001010: solve_cell = 0;
            9'b110001011: solve_cell = 0;
            9'b110001100: solve_cell = 0;
            9'b110001101: solve_cell = 0;
            9'b110001110: solve_cell = 0;
            9'b110001111: solve_cell = 0;
            9'b110010000: solve_cell = 1;
            9'b110010001: solve_cell = 1;
            9'b110010010: solve_cell = 1;
            9'b110010011: solve_cell = 0;
            9'b110010100: solve_cell = 1;
            9'b110010101: solve_cell = 0;
            9'b110010110: solve_cell = 0;
            9'b110010111: solve_cell = 0;
            9'b110011000: solve_cell = 1;
            9'b110011001: solve_cell = 0;
            9'b110011010: solve_cell = 0;
            9'b110011011: solve_cell = 0;
            9'b110011100: solve_cell = 0;
            9'b110011101: solve_cell = 0;
            9'b110011110: solve_cell = 0;
            9'b110011111: solve_cell = 0;
            9'b110100000: solve_cell = 1;
            9'b110100001: solve_cell = 0;
            9'b110100010: solve_cell = 0;
            9'b110100011: solve_cell = 0;
            9'b110100100: solve_cell = 0;
            9'b110100101: solve_cell = 0;
            9'b110100110: solve_cell = 0;
            9'b110100111: solve_cell = 0;
            9'b110101000: solve_cell = 0;
            9'b110101001: solve_cell = 0;
            9'b110101010: solve_cell = 0;
            9'b110101011: solve_cell = 0;
            9'b110101100: solve_cell = 0;
            9'b110101101: solve_cell = 0;
            9'b110101110: solve_cell = 0;
            9'b110101111: solve_cell = 0;
            9'b110110000: solve_cell = 1;
            9'b110110001: solve_cell = 0;
            9'b110110010: solve_cell = 0;
            9'b110110011: solve_cell = 0;
            9'b110110100: solve_cell = 0;
            9'b110110101: solve_cell = 0;
            9'b110110110: solve_cell = 0;
            9'b110110111: solve_cell = 0;
            9'b110111000: solve_cell = 0;
            9'b110111001: solve_cell = 0;
            9'b110111010: solve_cell = 0;
            9'b110111011: solve_cell = 0;
            9'b110111100: solve_cell = 0;
            9'b110111101: solve_cell = 0;
            9'b110111110: solve_cell = 0;
            9'b110111111: solve_cell = 0;
            9'b111000000: solve_cell = 1;
            9'b111000001: solve_cell = 0;
            9'b111000010: solve_cell = 0;
            9'b111000011: solve_cell = 0;
            9'b111000100: solve_cell = 0;
            9'b111000101: solve_cell = 0;
            9'b111000110: solve_cell = 0;
            9'b111000111: solve_cell = 0;
            9'b111001000: solve_cell = 0;
            9'b111001001: solve_cell = 0;
            9'b111001010: solve_cell = 0;
            9'b111001011: solve_cell = 0;
            9'b111001100: solve_cell = 0;
            9'b111001101: solve_cell = 0;
            9'b111001110: solve_cell = 0;
            9'b111001111: solve_cell = 0;
            9'b111010000: solve_cell = 1;
            9'b111010001: solve_cell = 0;
            9'b111010010: solve_cell = 0;
            9'b111010011: solve_cell = 0;
            9'b111010100: solve_cell = 0;
            9'b111010101: solve_cell = 0;
            9'b111010110: solve_cell = 0;
            9'b111010111: solve_cell = 0;
            9'b111011000: solve_cell = 0;
            9'b111011001: solve_cell = 0;
            9'b111011010: solve_cell = 0;
            9'b111011011: solve_cell = 0;
            9'b111011100: solve_cell = 0;
            9'b111011101: solve_cell = 0;
            9'b111011110: solve_cell = 0;
            9'b111011111: solve_cell = 0;
            9'b111100000: solve_cell = 0;
            9'b111100001: solve_cell = 0;
            9'b111100010: solve_cell = 0;
            9'b111100011: solve_cell = 0;
            9'b111100100: solve_cell = 0;
            9'b111100101: solve_cell = 0;
            9'b111100110: solve_cell = 0;
            9'b111100111: solve_cell = 0;
            9'b111101000: solve_cell = 0;
            9'b111101001: solve_cell = 0;
            9'b111101010: solve_cell = 0;
            9'b111101011: solve_cell = 0;
            9'b111101100: solve_cell = 0;
            9'b111101101: solve_cell = 0;
            9'b111101110: solve_cell = 0;
            9'b111101111: solve_cell = 0;
            9'b111110000: solve_cell = 0;
            9'b111110001: solve_cell = 0;
            9'b111110010: solve_cell = 0;
            9'b111110011: solve_cell = 0;
            9'b111110100: solve_cell = 0;
            9'b111110101: solve_cell = 0;
            9'b111110110: solve_cell = 0;
            9'b111110111: solve_cell = 0;
            9'b111111000: solve_cell = 0;
            9'b111111001: solve_cell = 0;
            9'b111111010: solve_cell = 0;
            9'b111111011: solve_cell = 0;
            9'b111111100: solve_cell = 0;
            9'b111111101: solve_cell = 0;
            9'b111111110: solve_cell = 0;
            9'b111111111: solve_cell = 0;
            default: solve_cell = 0;
        endcase;
    end
    endfunction;
    
    generate
    for (genvar i = 0; i <= map_width*(map_width - 1); i = i + map_width) begin
        for (genvar j = 0; j < map_width; j = j + 1) begin
            if (i + j == 0)
                assign next_state[i + j] = solve_cell({4'b0000, state[i + j], state[i + j + 1], 1'b0, state[i + j + map_width], state[i + j + map_width + 1]});
            else if (i == 0 && j > 0 && j < map_width - 1)
                assign next_state[i + j] = solve_cell({3'b000, state[i + j - 1], state[i + j], state[i + j + 1], state[i + j + map_width - 1], state[i + j + map_width], state[i + j + map_width + 1]});
            else if (i + j == map_width - 1)
                assign next_state[i + j] = solve_cell({3'b000, state[i + j - 1], state[i + j], 1'b0, state[i + j + map_width - 1], state[i + j + map_width], 1'b0});
            else if (i > 0 && i < map_width*(map_width - 1) && j == 0)
                assign next_state[i + j] = solve_cell({1'b0, state[i + j - map_width], state[i + j - map_width + 1], 1'b0, state[i + j], state[i + j + 1], 1'b0, state[i + j + map_width], state[i + j + map_width + 1]});
            else if (i > 0 && i < map_width*(map_width - 1) && j == map_width - 1)
                assign next_state[i + j] = solve_cell({state[i + j - map_width - 1], state[i + j - map_width], 1'b0, state[i + j - 1], state[i + j], 1'b0, state[i + j + map_width - 1], state[i + j + map_width], 1'b0});
            else if (i + j == map_width*(map_width - 1))
                assign next_state[i + j] = solve_cell({1'b0, state[i + j - map_width], state[i + j - map_width + 1], 1'b0, state[i + j], state[i + j + 1], 3'b000});
            else if (i == map_width*(map_width - 1) && j > 0 && j < map_width - 1)
                assign next_state[i + j] = solve_cell({state[i + j - map_width - 1], state[i + j - map_width], state[i + j - map_width + 1], state[i + j - 1], state[i + j], state[i + j + 1], 3'b000});
            else if (i + j == map_width*map_width - 1)
                assign next_state[i + j] = solve_cell({state[i + j - map_width - 1], state[i + j - map_width], 1'b0, state[i + j - 1], state[i + j], 1'b0, 3'b000});
            else
                assign next_state[i + j] = solve_cell({state[i + j - map_width - 1], state[i + j - map_width], state[i + j - map_width + 1], state[i + j - 1], state[i + j], state[i + j + 1], state[i + j + map_width - 1], state[i + j + map_width], state[i + j + map_width + 1]});
        end
    end
    endgenerate
    
endmodule
